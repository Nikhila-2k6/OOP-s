// Code your testbench here
// or browse Examples
//custom constructor is for memory creation
//if not using custom constructor we will create two handles which increases the complexity

class vlsi;
  int data; //class member /data member
  bit [7:0]data1;
  shortint data2;
  function new(input int datain=0,input bit [7:0]datain1=8'h00,input shortint datain2=0);
    data=datain; //class member=function custom constructor argument
    data1=datain1;
    data2=datain2;
  endfunction
endclass

module tb;
  vlsi v;
  initial begin
    v=new(31,20,19); //object creation / new is called constructor
    $display("data=%0d,data1=%0d,data2=%0d",v.data,v.data1,v.data2);
  end
endmodule
  //output:
# KERNEL: data=31,data1=20,data2=19
